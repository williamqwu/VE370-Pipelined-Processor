// pipelined register for ID/EX stage

`timescale 1ns / 1ps

module pr_id_ex(

);

endmodule
