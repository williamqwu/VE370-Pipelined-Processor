// pipelined register for MEM/WB stage

`timescale 1ns / 1ps

module pr_mem_wb(

);

endmodule
