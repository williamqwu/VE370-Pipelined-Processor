// main driver program for single-cycle processor

module main(
  input clk
);

  // TODO

endmodule
