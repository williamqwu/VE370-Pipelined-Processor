// pipelined register for EX/MEM stage

`timescale 1ns / 1ps

module pr_ex_mem(

);

endmodule
