// pipelined register for IF/ID stage

`timescale 1ns / 1ps

module pr_if_id(

);

endmodule
